// ----------------------------------------------------
// module regfile (Register file)
// ----------------------------------------------------

module regfile();

endmodule // 